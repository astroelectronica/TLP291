.title KiCad schematic
.include "C:/AE/TLP291/TLP291_SE.mod"
R1 0 /K {RK}
XU1 /IN /K 0 /OUT TLP291_SE
V1 /IN 0 PULSE( 0 {VPUL} {delay} {tr} {tf} {duty} {cycle} )
V2 VDD 0 DC {VSOURCE}
R2 /OUT VDD {RC}
.end
